`ifndef __OPCODE_VH__
`define __OPCODE_VH__

`define MOVI   4'b0000 
`define ADDI   4'b0001
`define ADD    4'b0010
`define SUB    4'b0011
`define ANDI   4'b0100
`define AND    4'b0101
`define OR     4'b0110
`define JUMP   4'b1000
`define LOAD   4'b1100
`define STORE  4'b1101

`endif

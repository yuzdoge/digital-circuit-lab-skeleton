`ifndef __ALUFUNC_VH__
`define __ALUFUNC_VH__

`define ALU_ADD     3'b000

`endif

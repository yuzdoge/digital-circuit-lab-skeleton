`ifndef __OPCODE_VH__
`define __OPCODE_VH__

`define MOVI 4'b0000 
`define MOVE 4'b0001
`define ADDI 4'b0010
`define ADD  4'b0011
`define SUB  4'b0101
`define ANDI 4'b0110
`define AND  4'b0111
`define OR   4'b1001
`define JUMP 4'b1010

`endif
